`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:26:49 12/02/2015 
// Design Name: 
// Module Name:    lab10
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab10(
  input clk,
  input reset,
  output [7:0] led,
  input ROT_A,
  input ROT_B,

  // VGA specific I/O ports
  output VGA_HSYNC,
  output VGA_VSYNC,
  output VGA_RED,
  output VGA_GREEN,
  output VGA_BLUE
  );
	
	localparam S_MAIN_WAIT = 0, S_MAIN_RESET = 1, S_MAIN_STORE = 2, S_MAIN_REPLACE = 3, S_MAIN_FINISH = 4, S_MAIN_CLEAR = 5;

  // Declare system variables
  reg [7:0] led_on[0:7];
  wire rot_event;
  wire rot_right;
	reg [2:0] pos;
	reg [16:0] addr_in;
	reg [16:0] addr_out;
	reg [12:0] counter_x;
	reg [12:0] counter_y;
	reg write;
	reg [15:0] clear;
	reg [12:0]tmp_counter;
	reg [12:0] x;
	reg [2:0]tmp[111:0];
	reg [3:0] P, P_next;
	reg [3:0]debug;
	integer i;

  // declare SRAM control signals
  wire [16:0] sram_addr;
  wire [2:0]  data_in;
  wire [2:0]  data_out;
  wire        we, en;

  // General VGA control signals
  wire video_on;      // when video_on is 0, the VGA controller is sending
                      // synchronization signals to the display device.

  wire pixel_tick;    // when pixel tick is 1, we must update the RGB value
                      // based for the new coordinate (pixel_x, pixel_y)

  wire [9:0] pixel_x; // x coordinate of the next pixel (between 0 ~ 639) 
  wire [9:0] pixel_y; // y coordinate of the next pixel (between 0 ~ 479)

  reg  [2:0] rgb_reg;  // RGB value for the current pixel
  reg  [2:0] rgb_next; // RGB value for the next pixel

  // Application-specific VGA signals
  reg  [16:0] dummy_addr;
  wire [2:0] current_rgb; // RGB values for the frame display application.
                          // In this demo, the value is generated by
                          // a video pattern generator:
                          //      video_pattern(id, x, y, current_rgb),
                          // where the input is the current scan coordinate (x, y),
                          // and the output is the RGB value of the video pattern
                          // 'id' at pixel (x, y).
  reg  [2:0] pattern_id;

  // Declare the video buffer size
  localparam VBUF_W = 320; // video buffer width
  localparam VBUF_H = 240; // video buffer height

  // Instiantiate a VGA sync signal generator
  vga_sync vs0(
    .clk(clk), .reset(reset), .oHS(VGA_HSYNC), .oVS(VGA_VSYNC),
    .visible(video_on), .p_tick(pixel_tick),
    .pixel_x(pixel_x), .pixel_y(pixel_y)
  );

  // Instiantiate a rotary dial controller
  Rotation_direction RTD(
    .CLK(clk),
    .ROT_A(ROT_A),
    .ROT_B(ROT_B),
    .rotary_event(rot_event),
    .rotary_right(rot_right)
  );

  // Instiantiate a video test pattern generator
  video_pattern vp0(
    .id(pattern_id),
    .x(pixel_x),
    .y(pixel_y),
    .rgb(current_rgb)
  );

  assign led = debug; // put data_out here to keep sram from being removed.

  // ------------------------------------------------------------------------
  // The following code describes an initialized SRAM memory block that
  // stores an 320x240 3-bit city image, plus a 112x40 moon image.
  sram #(.DATA_WIDTH(3), .ADDR_WIDTH(17), .RAM_SIZE(VBUF_W*VBUF_H+112*40))
    ram0 (.clk(clk), .we(we), .en(en),
            .addr(sram_addr), .data_i(data_in), .data_o(data_out));

  assign we = (P == S_MAIN_REPLACE || P == S_MAIN_CLEAR) ? 1 : 0; // SRAM is read-only for the sample code. You MUST change it for lab10.
  assign en = 1; // Always enable the SRAM block.
  assign sram_addr = (P == S_MAIN_WAIT) ? dummy_addr : ((P == S_MAIN_STORE) ? addr_out : addr_in);
  assign data_in = (P == S_MAIN_REPLACE) ? tmp[tmp_counter] : 3'b001; // SRAM is read-only so we tie inputs to zeros.
  // End of the SRAM memory block.
  // ------------------------------------------------------------------------
  always @ (posedge clk) begin
		if (reset)
		  dummy_addr <= 0;
		else if(P == S_MAIN_WAIT)
		  dummy_addr <= (pixel_x / 2) + (pixel_y / 2) * 320;
	end
	always@ (posedge clk) begin
		if(reset) P <= S_MAIN_CLEAR;////
		else P <= P_next;
	end
	
	always @(*) begin
		case(P) 
			S_MAIN_WAIT:
				if(rot_event)	P_next = S_MAIN_RESET;
				else if(reset)	P_next = S_MAIN_CLEAR;
				else P_next = S_MAIN_WAIT;
			S_MAIN_RESET:
				P_next = S_MAIN_STORE;
			S_MAIN_STORE:
				if(counter_x == 111) P_next = S_MAIN_REPLACE;
				else P_next = S_MAIN_STORE;
			S_MAIN_REPLACE:
				if(counter_y == 47) P_next = S_MAIN_FINISH;
				else if(tmp_counter == 111)P_next = S_MAIN_RESET;
				else P_next = S_MAIN_REPLACE;
			S_MAIN_FINISH:
				P_next = S_MAIN_WAIT;
			S_MAIN_CLEAR:
				if(clear == 320 * 48) P_next = S_MAIN_WAIT;
				else P_next = S_MAIN_CLEAR;
			default:P_next = S_MAIN_WAIT;
		endcase
	end
	
	always@ (posedge clk) begin
		if(reset) clear <= 0;
		else if(P == S_MAIN_CLEAR) begin
			debug <= 7;
			clear <= clear + 1;
		end
	end
	always@ (posedge clk) begin//////////addr_in/////////
		if(reset) addr_in <= 0;
		else if(P == S_MAIN_RESET) addr_in <= counter_y * 320 + pos * 32;
		else if(P == S_MAIN_REPLACE || P == S_MAIN_CLEAR) addr_in <= addr_in + 1;
	end
	
	always@ (posedge clk) begin//////////////addr_out/////////
		if(reset || P == S_MAIN_RESET) addr_out <= 320*240 + (counter_y - 8) * 112;
		else if(P == S_MAIN_STORE) addr_out <= addr_out + 1;
	end
	
	always@ (posedge clk) begin///////////tmp///////////
		if(P == S_MAIN_STORE) tmp[tmp_counter] <= data_out;
	end
	
	always@ (posedge clk) begin///////////counter_y///////////
		if(reset || P == S_MAIN_WAIT) counter_y <= 8;
		else if(counter_x == 111) counter_y <= counter_y + 1;
	end
	
	always@ (posedge clk) begin////////counter_x////////
		if(P == S_MAIN_RESET || P == S_MAIN_WAIT || counter_x == 111) counter_x <= 0;
		else if(P == S_MAIN_STORE) counter_x <= counter_x + 1;
	end
	
	always@ (posedge clk) begin/////////////tmp_counter////////
		if(tmp_counter == 111 || P == S_MAIN_RESET) tmp_counter <= 0;
		else if(P == S_MAIN_STORE) tmp_counter <= tmp_counter + 1;
		else if(P == S_MAIN_REPLACE) tmp_counter <= tmp_counter + 1;
	end
  // ------------------------------------------------------------------------
  // Use the rotary input to select the video pattern.
  always@ (posedge clk) begin
    if (reset)
      pattern_id <= 3'b000;
    else if (rot_event && !rot_right)
      pattern_id <= pattern_id + 1;
    else if (rot_event && rot_right)
      pattern_id <= pattern_id - 1;
  end
  // End of the rotary input code.
  // ------------------------------------------------------------------------

  // VGA color pixel generator
  assign {VGA_RED, VGA_GREEN, VGA_BLUE} = rgb_reg;

  always @(posedge clk) begin
    if (pixel_tick) rgb_reg <= rgb_next;
  end

  always @(*) begin
    if (~video_on)
      rgb_next = 3'b000; // Synchronization period, must set RGB values to zero.
    else
      rgb_next = data_out; // RGB value at (pixel_x, pixel_y)
  // End of the video data display code.
  // ------------------------------------------------------------------------
  end
		
	always@ (posedge clk) begin
    if (reset)
      pos <= 3'b000;
    else if (rot_event && rot_right && pos < 3'b111)
      pos <= pos + 1;
    else if (rot_event && !rot_right && pos > 3'b000)
      pos <= pos - 1;
  end

endmodule
